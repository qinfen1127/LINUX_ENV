//==========================================================================================================================
//  @File Name  :  tb.v
//  @File Type  :  verilog
//  @Author     :  Howard
//  @E-mail     :  qinfen1127@163.com
//  @Date       :  2024-07-03
//  @Function   :  
//==========================================================================================================================

//---------------------------------------------------------------------------------------------------------------------
// testbench file header
//---------------------------------------------------------------------------------------------------------------------
`timescale 1ns/1ps

module tb ;

endmodule

//---------------------------------------------------------------------------------------------------------------------
// 
//---------------------------------------------------------------------------------------------------------------------
