//======================================================================
// Copyright(c) 2020, Chengdu Sino Microelectronics Technology CO., LTD.
//                         All Right Reserved
//
// Created by     : hr_li
// Filename       : ram.v
// Created On     : 2020-04-28
// Last Modified  : 2020-04-28
//
// Description: 
//
// Version        Modified by        Date           Description
// 1              hr_li              2020-04-28     original
//
//======================================================================

module ram (/*autoarg*/
   // Outputs
   dout,
   // Inputs
   clk, wen, din, waddr, raddr
   );

//--------------------------------------------------------------------------------------------
//  parameter define
//--------------------------------------------------------------------------------------------
parameter					DWIDTH		=	8   		;
parameter					AWIDTH      =	10   		;

//--------------------------------------------------------------------------------------------
//  input & output
//--------------------------------------------------------------------------------------------
input						clk							;
input						wen							;
input  		[DWIDTH-1:0]	din							;
input  		[AWIDTH-1:0]	waddr						;
input  		[AWIDTH-1:0]	raddr						;

output 		[DWIDTH-1:0]	dout						;

//--------------------------------------------------------------------------------------------
//  reg define
//--------------------------------------------------------------------------------------------
reg			[DWIDTH-1:0]	ram			[2**AWIDTH-1:0] ;
reg			[AWIDTH-1:0]	raddr_reg					;

//--------------------------------------------------------------------------------------------
//  write operation
//--------------------------------------------------------------------------------------------
always@(posedge clk) begin
	if(wen) begin
		ram[waddr] <= din ;
	end
end

//--------------------------------------------------------------------------------------------
//  read operation
//--------------------------------------------------------------------------------------------
always@(posedge clk) begin
	raddr_reg <= raddr ;
end

assign  dout = ram[raddr_reg] ;

endmodule

